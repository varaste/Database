library ieee;
use ieee.std_logic_1164.all;
architecture behavior of unsigned1 is
begin
	q <= a + b;	--(2)
end;
