entity logical_alu is
port ( a,b : in  std_logic_vesactor(2 downto 0);
       alu_
