entity logical_alu is
port ( a,b : in  std_logic_vesactor(2 downto 0);
       alu_out: out std_logic_vector(3 downto 0));
end logical_alu;

architecture behav of logical_alu is
beg
       	   op="011" else
       	    
end behav;
