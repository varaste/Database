
begin
	q <= a + b;	--(2)
end;
